--VHDL code for Program counter
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pc_32 is
    port (
        clk : in std_logic;
        pc_in : in std_logic_vector(31 downto 0);
        pc_out : out std_logic_vector(31 downto 0)
    );
end pc_32;

architecture beh of pc_32 is
	
begin

    process (clk)
    begin
        
        if rising_edge(clk) then
    
            --if pc_in=(others=>"xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx") then
            --  pc_out<="00000000000000000000000000000000";
            --else
            --   pc_out<=pc_in;
            --end if;
            
            
            ---if pc_in/="00000000000000000000000000000000" then
              ----  pc_out <= pc_in;
              ----else
                ---pc_out <= "00000000000000000000000000000000";
              -----end if;
              
              
              
              
              case pc_in(31 downto 0) is 
              when "00000000000000000000000000000000" => pc_out <= "00000000000000000000000000000000";	
              when "00000000000000000000000000000100" => pc_out <= "00000000000000000000000000000100"; 
              when "00000000000000000000000000001000" => pc_out <= "00000000000000000000000000001000"; 
              when "00000000000000000000000000001100" => pc_out <= "00000000000000000000000000001100"; 
              when "00000000000000000000000000010000" => pc_out <= "00000000000000000000000000010000"; 
              when "00000000000000000000000000010100" => pc_out <= "00000000000000000000000000010100";	
              when "00000000000000000000000000011000" => pc_out <= "00000000000000000000000000011000";	
              when "00000000000000000000000000011100" => pc_out <= "00000000000000000000000000011100";	
              when "00000000000000000000000000100000" => pc_out <= "00000000000000000000000000100000";	
              when "00000000000000000000000000100100" => pc_out <= "00000000000000000000000000100100";	
              when "00000000000000000000000000101000" => pc_out <= "00000000000000000000000000101000";	
              
              when "00000000000000000000000010101100" => pc_out <= "00000000000000000000000010101100";	
              when "00000000000000000000000010110000" => pc_out <= "00000000000000000000000010110000";	
              when "00000000000000000000000010110100" => pc_out <= "00000000000000000000000010110100";	
              when "00000000000000000000000010111000" => pc_out <= "00000000000000000000000010111000";	
              when "00000000000000000000000010111100" => pc_out <= "00000000000000000000000010111100";	  
                 
                
                
              when others => pc_out <= (others => '0');  
              
              end case;
                            
               
              
              
              
              
              
              
              
            
            
        end if;
        
        
        
         
        
        
    end process;
        
            
end architecture beh;